//Divide 48MGHz into usable hertz for sound, play notes (boing? somehow)





module jumpAudio (
input logic clk,
output logic jumpSoundOut
);











endmodule 
