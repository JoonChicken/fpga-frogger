module text_gen (
    input  logic [7:0] char_addr,     // Character code (ASCII)
    input  logic [2:0] row_addr,      // Row within character (0-7)
    output logic [7:0] bitmap         // 8-bit bitmap for the row
);

    logic [7:0] rom [0:687];  // 256 chars * 8 rows = 2048 entries
    // 100 chars only in this rom bc no need for not alphanumeric
    
    initial begin
        // Initialize all characters to 0
        for (int i = 0; i < 687; i++) begin
            rom[i] = 8'b0;
        end
        
        // Define ANSI-style 8x8 font bitmaps
        
        // Space (ASCI - 32I 32)
        rom['h20*8 + 0 - 32] = 8'b00000000;
        rom['h20*8 + 1 - 32] = 8'b00000000;
        rom['h20*8 + 2 - 32] = 8'b00000000;
        rom['h20*8 + 3 - 32] = 8'b00000000;
        rom['h20*8 + 4 - 32] = 8'b00000000;
        rom['h20*8 + 5 - 32] = 8'b00000000;
        rom['h20*8 + 6 - 32] = 8'b00000000;
 
        // : (ASCII 58 - 32) - Colon
        rom['h3A*8 + 0 - 32] = 8'b00000000;  // 
        rom['h3A*8 + 1 - 32] = 8'b00110000;  //   ##
        rom['h3A*8 + 2 - 32] = 8'b00110000;  //   ##
        rom['h3A*8 + 3 - 32] = 8'b00000000;  // 
        rom['h3A*8 + 4 - 32] = 8'b00000000;  // 
        rom['h3A*8 + 5 - 32] = 8'b00110000;  //   ##
        rom['h3A*8 + 6 - 32] = 8'b00110000;  //   ##
 
        // 0 (ASCII 48 - 32)
        rom['h30*8 + 0 - 32] = 8'b01111000;  //  ####
        rom['h30*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h30*8 + 2 - 32] = 8'b11011100;  // ## ###
        rom['h30*8 + 3 - 32] = 8'b11111100;  // ######
        rom['h30*8 + 4 - 32] = 8'b11101100;  // ### ##
        rom['h30*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h30*8 + 6 - 32] = 8'b01111000;  //  ####
         
        // 1 (ASCII 49 - 32)
        rom['h31*8 + 0 - 32] = 8'b00110000;  //   ##
        rom['h31*8 + 1 - 32] = 8'b01110000;  //  ###
        rom['h31*8 + 2 - 32] = 8'b00110000;  //   ##
        rom['h31*8 + 3 - 32] = 8'b00110000;  //   ##
        rom['h31*8 + 4 - 32] = 8'b00110000;  //   ##
        rom['h31*8 + 5 - 32] = 8'b00110000;  //   ##
        rom['h31*8 + 6 - 32] = 8'b11111100;  // ######
         
        // 2 (ASCII 50 - 32)
        rom['h32*8 + 0 - 32] = 8'b01111000;  //  ####
        rom['h32*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h32*8 + 2 - 32] = 8'b00001100;  //     ##
        rom['h32*8 + 3 - 32] = 8'b00111000;  //   ###
        rom['h32*8 + 4 - 32] = 8'b01100000;  //  ##
        rom['h32*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h32*8 + 6 - 32] = 8'b11111100;  // ######
         
        // 3 (ASCII 51 - 32)
        rom['h33*8 + 0 - 32] = 8'b01111000;  //  ####
        rom['h33*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h33*8 + 2 - 32] = 8'b00001100;  //     ##
        rom['h33*8 + 3 - 32] = 8'b00111000;  //   ###
        rom['h33*8 + 4 - 32] = 8'b00001100;  //     ##
        rom['h33*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h33*8 + 6 - 32] = 8'b01111000;  //  ####
         
        // 4 (ASCII 52 - 32)
        rom['h34*8 + 0 - 32] = 8'b00011100;  //    ###
        rom['h34*8 + 1 - 32] = 8'b00111100;  //   ####
        rom['h34*8 + 2 - 32] = 8'b01101100;  //  ## ##
        rom['h34*8 + 3 - 32] = 8'b11001100;  // ##  ##
        rom['h34*8 + 4 - 32] = 8'b11111110;  // #######
        rom['h34*8 + 5 - 32] = 8'b00001100;  //     ##
        rom['h34*8 + 6 - 32] = 8'b00011110;  //    ####
         
        // 5 (ASCII 53 - 32)
        rom['h35*8 + 0 - 32] = 8'b11111100;  // ######
        rom['h35*8 + 1 - 32] = 8'b11000000;  // ##
        rom['h35*8 + 2 - 32] = 8'b11111000;  // #####
        rom['h35*8 + 3 - 32] = 8'b00001100;  //     ##
        rom['h35*8 + 4 - 32] = 8'b00001100;  //     ##
        rom['h35*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h35*8 + 6 - 32] = 8'b01111000;  //  ####
         
        // 6 (ASCII 54 - 32)
        rom['h36*8 + 0 - 32] = 8'b00111000;  //   ###
        rom['h36*8 + 1 - 32] = 8'b01100000;  //  ##
        rom['h36*8 + 2 - 32] = 8'b11000000;  // ##
        rom['h36*8 + 3 - 32] = 8'b11111000;  // #####
        rom['h36*8 + 4 - 32] = 8'b11001100;  // ##  ##
        rom['h36*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h36*8 + 6 - 32] = 8'b01111000;  //  ####
         
        // 7 (ASCII 55 - 32)
        rom['h37*8 + 0 - 32] = 8'b11111100;  // ######
        rom['h37*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h37*8 + 2 - 32] = 8'b00001100;  //     ##
        rom['h37*8 + 3 - 32] = 8'b00011000;  //    ##
        rom['h37*8 + 4 - 32] = 8'b00110000;  //   ##
        rom['h37*8 + 5 - 32] = 8'b00110000;  //   ##
        rom['h37*8 + 6 - 32] = 8'b00110000;  //   ##
         
        // 8 (ASCII 56 - 32)
        rom['h38*8 + 0 - 32] = 8'b01111000;  //  ####
        rom['h38*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h38*8 + 2 - 32] = 8'b11001100;  // ##  ##
        rom['h38*8 + 3 - 32] = 8'b01111000;  //  ####
        rom['h38*8 + 4 - 32] = 8'b11001100;  // ##  ##
        rom['h38*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h38*8 + 6 - 32] = 8'b01111000;  //  ####
         
        // 9 (ASCII 57 - 32)
        rom['h39*8 + 0 - 32] = 8'b01111000;  //  ####
        rom['h39*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h39*8 + 2 - 32] = 8'b11001100;  // ##  ##
        rom['h39*8 + 3 - 32] = 8'b01111100;  //  #####
        rom['h39*8 + 4 - 32] = 8'b00001100;  //     ##
        rom['h39*8 + 5 - 32] = 8'b00011000;  //    ##
        rom['h39*8 + 6 - 32] = 8'b01110000;  //  ###
     
        // F (ASCII 70 - 32)
        rom['h46*8 + 0 - 32] = 8'b11111100;  // ######
        rom['h46*8 + 1 - 32] = 8'b11000000;  // ##
        rom['h46*8 + 2 - 32] = 8'b11000000;  // ##
        rom['h46*8 + 3 - 32] = 8'b11111000;  // #####
        rom['h46*8 + 4 - 32] = 8'b11000000;  // ##
        rom['h46*8 + 5 - 32] = 8'b11000000;  // ##
        rom['h46*8 + 6 - 32] = 8'b11000000;  // ##
     
        // G (ASCII 71 - 32)
        rom['h47*8 + 0 - 32] = 8'b01111100;  //  #####
        rom['h47*8 + 1 - 32] = 8'b11000110;  // ##   ##
        rom['h47*8 + 2 - 32] = 8'b11000000;  // ##
        rom['h47*8 + 3 - 32] = 8'b11011110;  // ## ####
        rom['h47*8 + 4 - 32] = 8'b11000110;  // ##   ##
        rom['h47*8 + 5 - 32] = 8'b11000110;  // ##   ##
        rom['h47*8 + 6 - 32] = 8'b01111100;  //  #####
     
        rom['h48*8 + 0 - 32] = 8'b11001100;  // ##  ##
        rom['h48*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h48*8 + 2 - 32] = 8'b11001100;  // ##  ##
        rom['h48*8 + 3 - 32] = 8'b11111100;  // ######
        rom['h48*8 + 4 - 32] = 8'b11001100;  // ##  ##
        rom['h48*8 + 5 - 32] = 8'b11001100;  // ##  ##
        rom['h48*8 + 6 - 32] = 8'b11001100;  // ##  ##
     
        rom['h49*8 + 0 - 32] = 8'b11111100;  // ######
        rom['h49*8 + 1 - 32] = 8'b00110000;  //   ##
        rom['h49*8 + 2 - 32] = 8'b00110000;  //   ##
        rom['h49*8 + 3 - 32] = 8'b00110000;  //   ##
        rom['h49*8 + 4 - 32] = 8'b00110000;  //   ##
        rom['h49*8 + 5 - 32] = 8'b00110000;  //   ##
        rom['h49*8 + 6 - 32] = 8'b11111100;  // ######
 
        rom['h4C*8 + 0 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 1 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 2 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 3 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 4 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 5 - 32] = 8'b11000000;  // ##
        rom['h4C*8 + 6 - 32] = 8'b11111100;  // ######
 
        rom['h56*8 + 0 - 32] = 8'b11001100;  // ##  ##
        rom['h56*8 + 1 - 32] = 8'b11001100;  // ##  ##
        rom['h56*8 + 2 - 32] = 8'b11001100;  // ##  ##
        rom['h56*8 + 3 - 32] = 8'b11001100;  // ##  ##
        rom['h56*8 + 4 - 32] = 8'b11001100;  // ##  ##
        rom['h56*8 + 5 - 32] = 8'b01111000;  //  ####
        rom['h56*8 + 6 - 32] = 8'b00110000;  //   ##
         
        // P (ASCII 80 - 32)
        rom['h50*8 + 0 - 32] = 8'b11111000;
        rom['h50*8 + 1 - 32] = 8'b11001100;
        rom['h50*8 + 2 - 32] = 8'b11001100;
        rom['h50*8 + 3 - 32] = 8'b11111000;
        rom['h50*8 + 4 - 32] = 8'b11000000;
        rom['h50*8 + 5 - 32] = 8'b11000000;
        rom['h50*8 + 6 - 32] = 8'b11000000;
         
        // R (ASCII 82 - 32)
        rom['h52*8 + 0 - 32] = 8'b11111000;
        rom['h52*8 + 1 - 32] = 8'b11001100;
        rom['h52*8 + 2 - 32] = 8'b11001100;
        rom['h52*8 + 3 - 32] = 8'b11111000;
        rom['h52*8 + 4 - 32] = 8'b11011000;
        rom['h52*8 + 5 - 32] = 8'b11001100;
        rom['h52*8 + 6 - 32] = 8'b11000110;
         
        // E (ASCII 69 - 32)
        rom['h45*8 + 0 - 32] = 8'b11111100;
        rom['h45*8 + 1 - 32] = 8'b11000000;
        rom['h45*8 + 2 - 32] = 8'b11000000;
        rom['h45*8 + 3 - 32] = 8'b11111000;
        rom['h45*8 + 4 - 32] = 8'b11000000;
        rom['h45*8 + 5 - 32] = 8'b11000000;
        rom['h45*8 + 6 - 32] = 8'b11111100;
         
        // S (ASCII 83 - 32)
        rom['h53*8 + 0 - 32] = 8'b01111100;
        rom['h53*8 + 1 - 32] = 8'b11000110;
        rom['h53*8 + 2 - 32] = 8'b11000000;
        rom['h53*8 + 3 - 32] = 8'b01111100;
        rom['h53*8 + 4 - 32] = 8'b00000110;
        rom['h53*8 + 5 - 32] = 8'b11000110;
        rom['h53*8 + 6 - 32] = 8'b01111100;
         
        // A (ASCII 65 - 32)
        rom['h41*8 + 0 - 32] = 8'b00110000;
        rom['h41*8 + 1 - 32] = 8'b01111000;
        rom['h41*8 + 2 - 32] = 8'b11001100;
        rom['h41*8 + 3 - 32] = 8'b11001100;
        rom['h41*8 + 4 - 32] = 8'b11111100;
        rom['h41*8 + 5 - 32] = 8'b11001100;
        rom['h41*8 + 6 - 32] = 8'b11001100;
         
        // N (ASCII 78 - 32)
        rom['h4E*8 + 0 - 32] = 8'b11001100;
        rom['h4E*8 + 1 - 32] = 8'b11101100;
        rom['h4E*8 + 2 - 32] = 8'b11111100;
        rom['h4E*8 + 3 - 32] = 8'b11111100;
        rom['h4E*8 + 4 - 32] = 8'b11011100;
        rom['h4E*8 + 5 - 32] = 8'b11001100;
        rom['h4E*8 + 6 - 32] = 8'b11001100;
         
        // Y (ASCII 89 - 32)
        rom['h59*8 + 0 - 32] = 8'b11001100;
        rom['h59*8 + 1 - 32] = 8'b11001100;
        rom['h59*8 + 2 - 32] = 8'b11001100;
        rom['h59*8 + 3 - 32] = 8'b01111000;
        rom['h59*8 + 4 - 32] = 8'b00110000;
        rom['h59*8 + 5 - 32] = 8'b00110000;
        rom['h59*8 + 6 - 32] = 8'b00110000;
         
        // K (ASCII 75 - 32)
        rom['h4B*8 + 0 - 32] = 8'b11001100;
        rom['h4B*8 + 1 - 32] = 8'b11011000;
        rom['h4B*8 + 2 - 32] = 8'b11110000;
        rom['h4B*8 + 3 - 32] = 8'b11100000;
        rom['h4B*8 + 4 - 32] = 8'b11110000;
        rom['h4B*8 + 5 - 32] = 8'b11011000;
        rom['h4B*8 + 6 - 32] = 8'b11001100;
         
        // T (ASCII 84 - 32)
        rom['h54*8 + 0 - 32] = 8'b11111100;
        rom['h54*8 + 1 - 32] = 8'b00110000;
        rom['h54*8 + 2 - 32] = 8'b00110000;
        rom['h54*8 + 3 - 32] = 8'b00110000;
        rom['h54*8 + 4 - 32] = 8'b00110000;
        rom['h54*8 + 5 - 32] = 8'b00110000;
        rom['h54*8 + 6 - 32] = 8'b00110000;
         
        // O (ASCII 79 - 32)
        rom['h4F*8 + 0 - 32] = 8'b01111000;
        rom['h4F*8 + 1 - 32] = 8'b11001100;
        rom['h4F*8 + 2 - 32] = 8'b11001100;
        rom['h4F*8 + 3 - 32] = 8'b11001100;
        rom['h4F*8 + 4 - 32] = 8'b11001100;
        rom['h4F*8 + 5 - 32] = 8'b11001100;
        rom['h4F*8 + 6 - 32] = 8'b01111000;
        

    end
    
    // Read from ROM
    assign bitmap = rom[{char_addr -32, row_addr}];

endmodule