//Divide 48MGHz into usable hertz for sound, play notes (womp-womp?)






module loseAudio (
input logic clk,
output logic loseSoundOut
);











endmodule 
