//Divide 48MGHz into usable hertz for sound, play notes (ta-da?)





module winAudio (
    input logic enable,
    input logic clk,
    output logic winSoundOut
);











endmodule 